module normips (CLOCKAUTO,ENTER1, SWITCH, RESET,/* RESET, BOTAO, *//*SWITCH, ENDERECO_INSTRUCAO_TEST, INSTRUCAO_TEST, 
					 BANCOREG_CONTROL_TEST, MEMDADOS_CONTROL_TEST, 
					 MUX1_CONTROL_TEST, MUX2_CONTROL_TEST, MUX3_CONTROL_TEST,
					 SAIDA_MUX1_TEST, SAIDA_MUX3_TEST, SAIDA_RD_TEST,
					 SAIDA_RS_TEST, SAIDA_RT_TEST, EXTENDIDO_TEST,
					 SAIDA_MUX2_TEST, ALU_RESULT_TEST, ALU_CONTROL_TEST,
					 MEMDADOS_SAIDA_TEST, EXTENDIDO2_TEST, EXTENDIDO_DESLOCADO_TEST,
					 SAIDA_MUX4_TEST, MUX4_CONTROL_TEST*/ SAIDA_MEMDADOS_TEST, UNIDADE, DEZENA,
					 CENTENA, MILHAR, D_MILHAR, C_MILHAR, MILHAO, D_MILHAO, UNIDADE2, DEZENA2, CENTENA2, MILHAR2, D_MILHAR2, C_MILHAR2, MILHAO2, 
											D_MILHAO2, INSTRUCAO_TEST, SAIDA_MUX4_TEST, RESULTADO_ALU_TEST,
					 SAIDA_MUX2_TEST, SAIDA_MUXN_TEST, SAIDA_MUX3_TEST, SAIDA_D1_TEST, SAIDA_D2_TEST, ENDERECO_INSTRUCAO_TEST, SAIDA_SWR_TEST);
					 
	input CLOCKAUTO;//, RESET;
	input ENTER1;
	input [15:0] SWITCH;
	input RESET;

	wire ENTER;
	wire ENTER2;
	
	output reg [31:0] INSTRUCAO_TEST;
	output reg [31:0] RESULTADO_ALU_TEST;
	output reg [31:0] SAIDA_MEMDADOS_TEST;
	output reg [31:0] SAIDA_MUXN_TEST;
	output reg [31:0] SAIDA_MUX4_TEST;
	output reg [31:0] SAIDA_MUX3_TEST;
	output reg [31:0] SAIDA_MUX2_TEST;
	output reg [31:0] SAIDA_D1_TEST;
	output reg [31:0] SAIDA_D2_TEST;
	output reg [31:0] ENDERECO_INSTRUCAO_TEST;
	output reg [31:0] SAIDA_SWR_TEST;

	wire CLOCK;
	wire [31:0] SAIDA_MUX4;
	wire [31:0] SAIDA_MUX3;
	wire [31:0] SAIDA_MUX2;
	wire [31:0] SAIDA_MUXN;
	wire [31:0] ENDERECO_INSTRUCAO;
	wire [31:0] INSTRUCAO;
	wire [31:0] ENDERECO;
	wire [31:0] SAIDA_D1;
	wire [31:0] SAIDA_D2;
	wire [31:0] SAIDA_SWR;
	wire [31:0] EXTENDIDO;
	wire [31:0] ALU_RESULT;
	wire [31:0] SAIDA_MEMDADOS;
	wire [31:0] EXTENDIDO2;
	wire SINAL_ZERO;
	wire SINAL_NEG;
	wire [3:0] CONTROLE_ALU;
	wire [2:0] CONTROLE_MUX4;
	wire [1:0] CONTROLE_MUX3;
	wire [1:0] CONTROLE_MUXN;
	wire CONTROLE_MUX2;
	wire CONTROLE_ESCRITA_BR;
	wire CONTROLE_ESCRITA_MEMDADOS;
	wire CONTROLE_JAL;
	wire CONTROLE_D2;
	wire CONTROLE_OPT;
	wire HALT;

	output [6:0] UNIDADE, DEZENA, CENTENA, MILHAR, D_MILHAR, C_MILHAR, MILHAO, D_MILHAO;
	output [6:0] UNIDADE2, DEZENA2, CENTENA2, MILHAR2, D_MILHAR2, C_MILHAR2, MILHAO2, D_MILHAO2;
	
	//freq_cut freq_cut(CLOCKAUTO, CLOCK);
	
	//debouncer debouncer(CLOCKAUTO, ~ENTER1, ENTER);
	
	//DeBounce DeBounce(CLOCKAUTO, 1, ENTER1, ENTER);
	temporizador temporizador(CLOCKAUTO, CLOCK);
	
	//one_shot_button one_shot_button(CLOCKAUTO, ENTER2, ENTER);
	
	programCounter programCounter(SAIDA_MUX4, ENDERECO_INSTRUCAO, CLOCK, /*~RESET,*/ ~RESET, HALT);
	
	memoriaInstrucao memoriaInstrucao(ENDERECO_INSTRUCAO, INSTRUCAO, CLOCK, ENDERECO, CLOCKAUTO);

	unidadeControle unidadeControle(INSTRUCAO[31:26], CLOCK, CONTROLE_MUX4, CONTROLE_MUX3, /*CONTROLE_MUX6,*/
											  CONTROLE_MUXN, CONTROLE_ALU, CONTROLE_MUX2, CONTROLE_ESCRITA_BR,
											  CONTROLE_D2, CONTROLE_ESCRITA_MEMDADOS, CONTROLE_OPT, CONTROLE_JAL, HALT, ~ENTER1);
	
	bancoRegistradores bancoRegistradores(INSTRUCAO[25:21], INSTRUCAO[20:16], INSTRUCAO[15:11], SAIDA_MUX3, SAIDA_D1,
													  SAIDA_D2, SAIDA_SWR, CONTROLE_ESCRITA_BR, CONTROLE_D2, CONTROLE_JAL, CLOCK, CLOCKAUTO);
													  
	extensor16_32 extensor16_32(INSTRUCAO[15:0], EXTENDIDO);
	extensor16_32 extensor13_32_SWITCHES(SWITCH, SWITCH_EXTENDIDO);

	MUX_2 MUX_2(SAIDA_D2, EXTENDIDO, SAIDA_MUX2, CONTROLE_MUX2);
	
	ALU ALU(SAIDA_D1, SAIDA_MUX2, ALU_RESULT, CONTROLE_ALU, SINAL_ZERO, SINAL_NEG, CLOCKAUTO);
	
	MUX_N MUX_N(ENDERECO, SAIDA_SWR, SAIDA_D1, EXTENDIDO, SAIDA_MUXN, CONTROLE_MUXN);

	memoriaDados memoriaDados(ALU_RESULT, SAIDA_MUXN, SAIDA_MEMDADOS, CONTROLE_ESCRITA_MEMDADOS, CLOCK, CLOCKAUTO);

	MUX_3 MUX_3(SAIDA_MEMDADOS, ALU_RESULT, EXTENDIDO, SWITCH_EXTENDIDO,SAIDA_MUX3, CONTROLE_MUX3);
	
	extensor26_28 extensor26_28(INSTRUCAO[25:0], EXTENDIDO2);
	
	MUX_4 MUX_4(ENDERECO_INSTRUCAO, EXTENDIDO, EXTENDIDO2, SAIDA_SWR, SAIDA_MUX4, CONTROLE_MUX4, SINAL_ZERO);
	
	output_normips output_normips(SAIDA_SWR, UNIDADE, DEZENA, CENTENA, MILHAR, D_MILHAR, C_MILHAR, MILHAO, 
											D_MILHAO, CLOCK, CONTROLE_OPT);
										
	output_normips output_normips2(ENDERECO_INSTRUCAO, UNIDADE2, DEZENA2, CENTENA2, MILHAR2, D_MILHAR2, C_MILHAR2, MILHAO2, 
											D_MILHAO2, CLOCK, 1'b1);
	
	always @ (posedge CLOCKAUTO) begin
		ENDERECO_INSTRUCAO_TEST = ENDERECO_INSTRUCAO;
		INSTRUCAO_TEST = INSTRUCAO;
		SAIDA_MEMDADOS_TEST = SAIDA_MEMDADOS;
		RESULTADO_ALU_TEST = ALU_RESULT;
		SAIDA_MUX4_TEST = SAIDA_MUX4;
		SAIDA_MUX2_TEST = SAIDA_MUX2;
		SAIDA_MUXN_TEST = SAIDA_MUXN;
		SAIDA_D1_TEST = SAIDA_D1;
		SAIDA_D2_TEST = SAIDA_D2;
		SAIDA_MUX3_TEST = SAIDA_MUX3;
		SAIDA_SWR_TEST = SAIDA_SWR;
	end
	
	
	
endmodule 