module jorgecore (CLOCK1, BTN, RESET, BOTAO, SWITCH, /*ENDERECO_INSTRUCAO_TEST, INSTRUCAO_TEST, 
					 BANCOREG_CONTROL_TEST, MEMDADOS_CONTROL_TEST, 
					 MUX1_CONTROL_TEST, MUX2_CONTROL_TEST, MUX3_CONTROL_TEST,
					 SAIDA_MUX1_TEST, SAIDA_MUX3_TEST, SAIDA_RD_TEST,
					 SAIDA_RS_TEST, SAIDA_RT_TEST, EXTENDIDO_TEST,
					 SAIDA_MUX2_TEST, ALU_RESULT_TEST, ALU_CONTROL_TEST,
					 MEMDADOS_SAIDA_TEST, EXTENDIDO2_TEST, EXTENDIDO_DESLOCADO_TEST,
					 SAIDA_MUX4_TEST, MUX4_CONTROL_TEST*/,UNIDADE, DEZENA,
					 CENTENA, MILHAR, D_MILHAR, C_MILHAR, MILHAO, D_MILHAO);
					 
	input CLOCK1, RESET;
	input BTN;
	input [15:0] SWITCH;
	input BOTAO;
	
	//wire CLOCK;
	wire [31:0] ENDERECO_INSTRUCAO;
	wire [31:0] INSTRUCAO;
	wire BANCOREG_CONTROL, MEMDADOS_CONTROL, MUX1_CONTROL, MUX2_CONTROL, SINAL_ZERO, SINAL_NEG;
	wire [1:0] MUX3_CONTROL;
	wire [4:0] SAIDA_MUX1;
	wire [31:0] SAIDA_MUX3;
	wire [31:0] SAIDA_RD;
	wire [31:0] SAIDA_RS;
	wire [31:0] SAIDA_RT;
	wire [31:0] EXTENDIDO;
	wire [31:0] SAIDA_MUX2;
	wire [31:0] ALU_RESULT;
	wire [2:0] ALU_CONTROL;
	wire [31:0] MEMDADOS_SAIDA;
	wire [31:0] EXTENDIDO2;
	wire [31:0] EXTENDIDO_DESLOCADO;
	wire [31:0] SAIDA_MUX4;
	wire [1:0] MUX4_CONTROL;
	wire HALT;
	wire MUX6_CONTROL;
	wire [15:0] SAIDA_MUX6;
	wire OPT_CONTROL;
	wire [31:0] SAIDA_MUX7;
	/*
	output [31:0] ENDERECO_INSTRUCAO_TEST;
	output [31:0] INSTRUCAO_TEST;
	output BANCOREG_CONTROL_TEST, MEMDADOS_CONTROL_TEST, MUX1_CONTROL_TEST, MUX2_CONTROL_TEST, MUX3_CONTROL_TEST;
	output [4:0] SAIDA_MUX1_TEST;
	output [31:0] SAIDA_MUX3_TEST;
	output [31:0] SAIDA_RD_TEST;
	output [31:0] SAIDA_RS_TEST;
	output [31:0] SAIDA_RT_TEST;
	output [31:0] EXTENDIDO_TEST;
	output [31:0] SAIDA_MUX2_TEST;
	output [31:0] ALU_RESULT_TEST;
	output [2:0] ALU_CONTROL_TEST;
	output [31:0] MEMDADOS_SAIDA_TEST;
	output [31:0] EXTENDIDO2_TEST;
	output [31:0] EXTENDIDO_DESLOCADO_TEST;
	output [31:0] SAIDA_MUX4_TEST;
	output [1:0] MUX4_CONTROL_TEST;
	*/
	output [6:0] UNIDADE, DEZENA, CENTENA, MILHAR, D_MILHAR, C_MILHAR, MILHAO, D_MILHAO;
	
	debouncer debouncer(CLOCK1, ~BTN, CLOCK);
	
	programCounter programCounter(SAIDA_MUX4, ENDERECO_INSTRUCAO, CLOCK, ~RESET, HALT);
	
	memoriaInstrucao memoriaInstrucao(ENDERECO_INSTRUCAO, INSTRUCAO, CLOCK);
	
	unidadeControle unidadeControle(INSTRUCAO[31:26], ~BOTAO, CLOCK, BANCOREG_CONTROL, MEMDADOS_CONTROL, 
											  MUX1_CONTROL, MUX2_CONTROL, MUX3_CONTROL, MUX4_CONTROL,
											  ALU_CONTROL, HALT, MUX6_CONTROL, OPT_CONTROL);
											  
	MUX_1 MUX_1(INSTRUCAO[20:16], INSTRUCAO[15:11], SAIDA_MUX1, MUX1_CONTROL);
	
	bancoRegistradores bancoRegistradores(INSTRUCAO[25:21], INSTRUCAO[20:16], SAIDA_MUX1, SAIDA_MUX3,
													  SAIDA_RD, SAIDA_RS, SAIDA_RT, BANCOREG_CONTROL, CLOCK);
													  
	MUX_6 MUX_6(INSTRUCAO[15:0], SWITCH, SAIDA_MUX6, MUX6_CONTROL);
	
	extensor16_32 extensor16_32(SAIDA_MUX6, EXTENDIDO);
	
	MUX_2 MUX_2(SAIDA_RT, EXTENDIDO, SAIDA_MUX2, MUX2_CONTROL);
	
	ALU ALU(SAIDA_RS, SAIDA_MUX2, ALU_RESULT, ALU_CONTROL, SINAL_ZERO, SINAL_NEG);
	
	memoriaDados memoriaDados(EXTENDIDO, SAIDA_RT, MEMDADOS_SAIDA, MEMDADOS_CONTROL, CLOCK);
	
	MUX_3 MUX_3(MEMDADOS_SAIDA, ALU_RESULT, EXTENDIDO, SAIDA_MUX3, MUX3_CONTROL);
	
	extensor26_28 extensor26_28(INSTRUCAO[25:0], EXTENDIDO2);
	
	MUX_4 MUX_4(ENDERECO_INSTRUCAO, EXTENDIDO, EXTENDIDO2, SAIDA_MUX4, MUX4_CONTROL, SINAL_ZERO);
	
	output_normips output_normips(SAIDA_RT, UNIDADE, DEZENA, CENTENA, MILHAR, D_MILHAR, C_MILHAR, MILHAO, 
											D_MILHAO, CLOCK, OPT_CONTROL);
	
	/*
	assign ENDERECO_INSTRUCAO_TEST = ENDERECO_INSTRUCAO;
	*/assign INSTRUCAO_TEST = INSTRUCAO;/*
	assign BANCOREG_CONTROL_TEST = BANCOREG_CONTROL;
	assign MEMDADOS_CONTROL_TEST = MEMDADOS_CONTROL;
	assign MUX1_CONTROL_TEST = MUX1_CONTROL;
	assign MUX2_CONTROL_TEST = MUX2_CONTROL;
	assign MUX3_CONTROL_TEST = MUX3_CONTROL;
	assign SAIDA_MUX1_TEST = SAIDA_MUX1;
	assign SAIDA_MUX3_TEST = SAIDA_MUX3;
	assign SAIDA_RD_TEST = SAIDA_RD;
	assign SAIDA_RS_TEST = SAIDA_RS;
	assign SAIDA_RT_TEST = SAIDA_RT;
	assign EXTENDIDO_TEST = EXTENDIDO;
	assign SAIDA_MUX2_TEST = SAIDA_MUX2;
	assign ALU_RESULT_TEST = ALU_RESULT;
	assign ALU_CONTROL_TEST = ALU_CONTROL;
	assign MEMDADOS_SAIDA_TEST = MEMDADOS_SAIDA;
	assign EXTENDIDO2_TEST = EXTENDIDO2;
	assign EXTENDIDO_DESLOCADO_TEST = EXTENDIDO_DESLOCADO;
	assign SAIDA_MUX4_TEST = SAIDA_MUX4;
	assign MUX4_CONTROL_TEST = MUX4_CONTROL;
	*/
endmodule 